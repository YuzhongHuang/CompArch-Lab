module finitestatemachine 
(
	input cs;
	input sclk;
	input rw;
);