module concat
(
	input[3:0] PC,
	input[25:0] dout,
	input[1:0] b00
);

